library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity q1 is
  port (
	X,Y,Z : in  STD_LOGIC;
	A : out STD_LOGIC := '0'	);
end entity;

architecture  rtl OF q1 IS

begin

end architecture;
