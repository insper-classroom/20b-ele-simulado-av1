library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity q2 is
  port (
    x    : in  STD_LOGIC_VECTOR(1 downto 0);
    y    : in  STD_LOGIC_VECTOR(1 downto 0);
    xeqy : out STD_LOGIC;
    xlty : out STD_LOGIC);
end entity;

architecture  rtl OF q2 IS

begin


end architecture;
